module Cont_M10(input logic clk, rst,
					 output logic [3:0] cont);

					 

	always@(posedge clk)
		begin
		
		end

endmodule
