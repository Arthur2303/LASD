`include "RegisterFile.sv"

module tb_ RegisterFile();

    // Inputs
    logic [N-1:0] wd3;
    logic [2:0] wa3, ra1, ra2;
    logic we3, clk, rst;
    //Outputs
    logic [N-1:0] rd1, rd2;





endmodule