module InstrMemory(	input logic  [7:0]   A,
							output logic [31:0] RD);
							
	always_comb
		begin
			case (A)
				8'b00000000: RD = 32'b001000_00000_00001_00000_00000_000011; // ADDi $1, $0, 3
				8'b00000001: RD = 32'b001000_00000_00010_00000_00000_001001; // ADDi $2, $0, 9
				8'b00000010: RD = 32'b000101_00001_00010_00000_00000_000010; // BNE $2, $1, 2
				8'b00000011: RD = 32'b000000_00001_00010_00011_00000_100100; // AND $3, $1, $2
				8'b00000100: RD = 32'b000000_00001_00010_00100_00000_100101; // OR $4, $1, $2
				8'b00000101: RD = 32'b000000_00001_00010_00101_00000_100111; // NOR $5, $1, $2
				8'b00000110: RD = 32'b000000_00101_00100_00110_00000_101010; // SLT $6, $5, $4
				8'b00001000: RD = 32'b001000_00000_00110_00000_00000_000101; // ADDi $6, $0, 5
				default: 	 RD = 32'b001000_00000_00111_00000_00000_000111; // ADDi $7, $0, 7 
			endcase	
		end
	
endmodule
