library verilog;
use verilog.vl_types.all;
entity tb_RegisterFile is
end tb_RegisterFile;
