module desafio();


endmodule
